library verilog;
use verilog.vl_types.all;
entity instr_register_test is
end instr_register_test;
